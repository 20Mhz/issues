module test (clk, in, out);
input clk;
input in;
output out;

  sky130_fd_sc_hd__dfxtp_4 _22045_ (
    .CLK(clk),
    .D(in),
    .Q(out )
  );
endmodule
